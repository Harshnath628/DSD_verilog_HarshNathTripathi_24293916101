`timescale 1ns / 1ps


module not_gate(
input a,
output res
    );
    assign res=~(a);
endmodule