`timescale 1ns / 1ps


module and_gate(
input a,b,
output res
    );
    assign res=(a&b);
endmodule