`timescale 1ns / 1ps


module tb_and(

    );
    reg a,b;
    wire res;
    and_gate uut(a,b,res);
    initial begin
    a=0;b=0;
    #10
    a=0;b=1;
    #10
    a=1;b=0;
    #10
    a=1;b=1;
    #10
    $finish;
    end
endmodule
